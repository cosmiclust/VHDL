library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity test_or_beh is
  Port ( a: in STD_LOGIC;
         b: in STD_LOGIC;
         c: in STD_LOGIC);
  end test_or_beh

architecture 
